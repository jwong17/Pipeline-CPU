`timescale 1ns / 1ps
`include "define.v"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:59:37 04/08/2016 
// Design Name: 
// Module Name:    dmemory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module dmemory(clk, rst, memwrite, memread, addr, data_in, fileid, data_out
    );
input clk;
  input rst;
  input memwrite;
  input memread;
  input [`ISIZE-1:0] addr;      // address input is 16 bit wide 
  input [`DSIZE-1:0] data_in;          // data input
  input [2:0] fileid;//file id selects which amoung the files given below (0-7 for different inputs for imem) and (8-16 for differnt D-mem inputs) for this lab we are using fileid=0
  output [`DSIZE-1:0] data_out;    // data output

  reg [`DSIZE-1:0] memory [0:32*`ISIZE-1]; //size of the memory
  reg [8*`MAX_LINE_LENGTH:0] line; /* Line of text read from file */

integer fin, i, c, r;
reg [`ISIZE-1:0] t_addr;
reg [`DSIZE-1:0] t_data;

reg [`ISIZE-1:0] addr_r;

assign data_out = memread ? memory[addr_r]: 16'b0;//Reading from the memory. Do note that there is a clock cycle delay for reading from the memory just to indicate that memories are slower.

  always @(posedge clk)
    begin
      if(rst)
        begin
	   addr_r <=0;
  	   case(fileid)
	        1: fin = $fopen("dmem_test0.txt","r");
        	2: fin = $fopen("dmem_test1.txt","r");
	        3: fin = $fopen("dmem_test2.txt","r");
        	4: fin = $fopen("dmem_test3.txt","r");
	        5: fin = $fopen("dmem_test4.txt","r");
        	6: fin = $fopen("dmem_test5.txt","r");
	        7: fin = $fopen("dmem_test6.txt","r");
		   8: fin = $fopen("dmem_test7.txt","r");
	  endcase
	  $write("Opening Fileid %d\n", fileid);

	  while(!$feof(fin)) begin
              c = $fgetc(fin);
              // check for comment
              if (c == "/" | c == "#" | c == "%")
                  r = $fgets(line, fin);
              else
                 begin
                    // Push the character back to the file then read the next time
                    r = $ungetc(c, fin);
                    r = $fscanf(fin, "%h %h",t_addr, t_data);
                    memory[t_addr]=t_data;
                 end
            end
            $fclose(fin);
	end
      else
        begin
	  addr_r <= addr;
          if (memwrite)// active-high write enable
            begin            
              memory[addr] <= data_in;
            end
	end
    end


endmodule
